module AMC1303Mx #(
    parameter SYSCLK_FREQ = 100_000_000
) (
    input logic resetn,    // active low reset, need to invert because
                           // dec256sinc24b is active high reset
    input logic sdat,
    
    output logic [15:0] out_data,
    output logic sclk
);

`timescale 1ns/1ps

//===================================================================
// Parameters and regs
//===================================================================
    localparam clk_period = 1000;    // 20MHz, 1000ns
    
    reg sysclk;    // clock generated by the ADC, 20MHz
    reg rst;       // inverted reset signal for the decimation filter
    reg [15:0] adcDat;    // connects the output of decimation filter 
                          // FIFO
                          
    reg [15:0] cdc1;      // output of first register in FIFO

//===================================================================
// Signal Assignment
//===================================================================    
assign rst = ~resetn;    // inverts the input reset low into a reset
                         // high the decimation filter uses

//===================================================================
// Architecture
//===================================================================

//===================================================================
// Decimation Filter
//===================================================================
dec256sinc24b #(
    .SYSCLK_FREQ(SYSCLK_FREQ)
) decimator (
    .mclk1(sclk),
    .reset(rst),
    .mdata1(sdat),
    .DATA(adcDat)
);

//===================================================================
// FIFO: 2 flipflops
//===================================================================
always_ff @( posedge sysclk ) begin : CDC
    cdc1 <= adcDat;
    out_data <= cdc1;    // output
end

//===================================================================
// clock generator
//===================================================================
initial sclk <= 0;
always #(clk_period/2) sclk <= ~sclk;

endmodule