//////////////////////////////////////////////////////////////////////////////////
// Company: RIT SPEX
// Engineer: Alexander Olds
// 
// Create Date: 03/29/2021 10:07:42 PM
// Design Name: 
// Module Name: LSM9DS1
// Project Name: urc_rover
// Target Devices: Artix 7 35T
// Tool Versions: Vivado 2020.2
// Description: LSM9DS1 IMU Driver & interpreter
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module LSM9DS1 #(
    parameter SYSCLK_FREQ = 100_000_000
) (
    input sclk,
    input rstn
);
    
endmodule